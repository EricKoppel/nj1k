title=NJ1K.org - Bestig New Jersey''s 52 berg över tusen fot
welcome.header=Välkommen!
welcometext=The New Jersey 1K Club is a fledgling organization that seeks to bring attention to the many hiking opportunities and challenges that the Garden State offers. New Hampshire has the AMC 4000''ers; the Adirondacks has its 46''ers; the Catskills and its 3500 Club. And now . . . New Jersey''s own peakbagging club: the 1K''ers. Sure, New Jersey''s great if you like diners, traffic, and an ever-entertaining political system, but don''t you ever have mountain envy? Ever wish you could climb a mountain around here and enjoy the progression of biomes? Ever wish you could break out the crampons and ice axe on Garden State mountains without worrying about wounding them? Ever wish you could have one of those cool peakbagger decals for New Jersey mountains like they have in our more vertically blessed states? Well, there''s nothing we can do to make New Jersey''s mountains any higher, and we don''t have the decals yet, but at the least we can have a New Jersey peakbagging club. Yeah, our mountains are less than lofty, but we''ve got a lot of them and a surprising number don''t even have trails to the tops.
copyright=Copyright © 2008-2013 Eric Koppel
most.recent.climbs=Senaste bestigningar
headlines=Nyheter
unknown=okänt

mountain.elevation=Höjd
mountain.decimal_degrees=Decimalgrader
mountain.county=County
mountain.ownership=Ägande
mountain.owner=Ägare
mountain.trail_map=Karta
mountain.topo=Topografisk karta
mountain.nhn=Nearest higher neighbor
mountain.others=Ascents of {0}
mountain.stats=Statistik
mountain.pictures.from=Bilder av {0}

ascent.title=Ascent of {0} ({2} feet) by {1}
ascent.trip_report=Trip report
ascent.pictures=Bilder
ascent.summit=Bergstopp
ascent.climber=Bestigare
ascent.mountain=Berg
ascent.date=Bestigningsdatum
ascent.successful=Successful
ascent.log=Log ascent
ascent.report=Trip report
ascent.pics=Ladda upp bilder
ascent.edit=Ändra ascent
ascent.climb.list=Bestigningslista
ascent.delete=Radera bestigning
ascent.delete.prompt=Are you sure you want to delete this ascent?

user.totalclimbs=Totala bestigningar
user.uniquesuccess=Unika bestigningar
user.percentcomplete=Procent klar

users.aspirants=Aspiranter

news.title=Rubrik
news.entry=Story
news.pics=Ladda upp bilder
news.edit=Redigera artikel
news.delete=Radera artikel
news.delete.prompt=Are you sure you want to delete this article?
news.date=Datum
news.nynjtc=Nyheter från NYNJTC

radius.title=Berg nära {0}
radius.search=Radius search
true=Ja
false=Nej

menu.news=Nyheter
menu.list=Listan
menu.members=Medlemmar
menu.links=Länkar
menu.login=Logga in
menu.logout=Logga ut
menu.register=Registrera
menu.news.submit=Submit News
menu.edit.account=Ditt konto
menu.ascent=Log Ascent
menu.contact=Kontakt
menu.about=Om oss

validation.email=This e-mail address is not registered
validation.email.taken=This e-mail address is already registered
validation.login.invalid=Ogiltig användarnamn eller lösenord
validation.passwords.equal=Passwords must match
validation.antispam=Not the highest point in New Jersey!

email=E-postadress
email.address=Din e-postadress
email.subject=Ämne
email.message=Meddelande
email.antispam=Anti-spam fråga. Vad heter New Jerseys högsta berg?
email.send=Skicka
email.sent=Tack för förfrågan!

name=Namn
password=Lösenord
password.reset=Begär nyttlösenord
password.forgot=Glömt lösenord?
confirmpassword=Bekräfta lösenord
aboutme=Om mig
profile.pic=Profilbild
account.updated=Ditt konto har uppdaterats

registration.success=Välkommen, {0}! You may now sign in.

welcome=Välkommen, {0}!

help.ascent.date=Ange bestigningsdatumet ({0}). Lämna tomt om datumet är okänt.
help.ascent.success=Did you make it to the top?
button.submit.ascent=Submit ascent
button.submit.login=Logga in
button.submit.news=Submit news

password.length=Lösenordet måste innehålla mellan 6 och 32 tecken
password.sent=Your new password has been sent to your e-mail address
mail.resetpassword.subject=Password reset
mail.resetpassword=You or someone has requested a password reset for your account on NJ1K.org. If you did not make this request, ignore this mail. Otherwise, log in with this temporary password: {0}
mail.message=You have received a message from {0}:\n\n{1}
cancel=Cancel
contact=Kontakta NJ1K Club
yes=Ja
no=Nej
about=Om